module seg7 #(parameter DELAY_RISE = 1, DELAY_FALL = 1)
(
    input [3:0] D,
    output reg [6:0] Q
);

always @(*)
begin
    case (D)
        4'b0000 : Q <= 7'b0111111; // 0
        4'b0001 : Q <= 7'b0000110; // 1
        4'b0010 : Q <= 7'b1011011; // 2
        4'b0011 : Q <= 7'b1001111; // 3
        4'b0100 : Q <= 7'b1100110; // 4
        4'b0101 : Q <= 7'b1101101; // 5
        4'b0110 : Q <= 7'b1111101; // 6
        4'b0111 : Q <= 7'b0000111; // 7
        4'b1000 : Q <= 7'b1111111; // 8
        4'b1001 : Q <= 7'b1101111; // 9

        // 4'b1010 : Q <= 7'b1110111; // A 
        // 4'b1011 : Q <= 7'b1111100; // B
        // 4'b1100 : Q <= 7'b1111001; // C
        // 4'b1101 : Q <= 7'10111110; // D
        // 4'b1110 : Q <= 7'b1111001; // E
        // 4'b1111 : Q <= 7'b1110001; // F
        
        default : Q <= 7'b1000000; // -
    endcase
end
endmodule

/*
        gfedcba
Q <= 7'b0000000;

  * * A * *
*           *
*           *
F           B
*           *
*           *
  * * G * * 
*           *
*           *
E           C
*           *
*           *
  * * D * *    *(DP)
DP not implemented
*/
